LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

PACKAGE tipos IS
  TYPE LOGIC_ARRAY_24_T IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR(23 downto 0);
  TYPE LOGIC_ARRAY_48_T IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR(47 downto 0);
  CONSTANT pa_k : integer := 3;
END tipos;
